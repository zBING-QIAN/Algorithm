library verilog;
use verilog.vl_types.all;
entity conv_if is
    port(
        clk             : in     vl_logic
    );
end conv_if;
