library verilog;
use verilog.vl_types.all;
entity mytb_sv_unit is
end mytb_sv_unit;
