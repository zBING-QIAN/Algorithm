library verilog;
use verilog.vl_types.all;
entity ntt_if is
    port(
        clk             : in     vl_logic;
        rst             : in     vl_logic
    );
end ntt_if;
